`define UART0_CLK_CTRL     8'h00
`define UART0_CTRL         8'h01
`define UART0_BAUD         8'h02
`define RST_FIFO0          8'h03
`define TX_FIFO0           8'h04
`define RX_FIFO0           8'h05
`define FIFO0_SZE          8'h06
`define FIFO0_STATUS       8'h07


`define GPIO_CTRL          8'h20
`define GPIO_OUT           8'h21
`define GPIO_STATUS        8'h22

`define MTIMECMP           8'h10
`define MCOUNTSTAR         8'h11 

`define SDStartAddr        8'h08
`define SDCounts           8'h09
`define DestAddr           8'h0a
`define DMAEN              8'h0b






